library verilog;
use verilog.vl_types.all;
entity tb_regC is
end tb_regC;
