library verilog;
use verilog.vl_types.all;
entity tb_instmem is
end tb_instmem;
