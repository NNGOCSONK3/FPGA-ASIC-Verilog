library verilog;
use verilog.vl_types.all;
entity tb_datamem is
end tb_datamem;
