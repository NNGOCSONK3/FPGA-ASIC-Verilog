library verilog;
use verilog.vl_types.all;
entity tb_PC is
end tb_PC;
