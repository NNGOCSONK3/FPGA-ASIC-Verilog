library verilog;
use verilog.vl_types.all;
entity tb_regA is
end tb_regA;
