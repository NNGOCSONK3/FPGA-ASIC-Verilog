library verilog;
use verilog.vl_types.all;
entity tb_regB is
end tb_regB;
